module PC (clock, in, out, LdPC, reset);
	input clock;
	input [15:0] in;
	output [15:0] out;
	
	

endmodule
